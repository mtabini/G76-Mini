parameter CLOCK_PHASE_SET_PIXEL_1     = 0;
parameter CLOCK_PHASE_READ_PIXEL_1    = 1;

parameter CLOCK_PHASE_SET_PIXEL_2     = 2;
parameter CLOCK_PHASE_READ_PIXEL_2    = 3;

parameter CLOCK_PHASE_READY_WRITE     = 4;
parameter CLOCK_PHASE_START_WRITE     = 5;

parameter CLOCK_PHASE_COMPLETE_WRITE  = 6;
parameter CLOCK_PHASE_IDLE_2          = 7;

parameter CLOCK_PHASE_RENDER_PIXEL_1  = 2;
parameter CLOCK_PHASE_RENDER_PIXEL_2  = 6;
