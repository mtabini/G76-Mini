  parameter
    CLOCK_PHASE_IDLE                = 0,
    CLOCK_PHASE_VIDEO_READ          = 1,
    CLOCK_PHASE_MEM_READ            = 2,
    CLOCK_PHASE_MEM_WRITE           = 3,
    CLOCK_PHASE_NOP                 = 4,
    CLOCK_PHASE_COMPLETE            = 5,

    CLOCK_PHASE_PREP_VIDEO_READ     = CLOCK_PHASE_COMPLETE,
    CLOCK_PHASE_PREP_MEMORY_OP      = CLOCK_PHASE_IDLE,
    CLOCK_PHASE_CLEAR_MEMORY_OP     = CLOCK_PHASE_COMPLETE;
